entity step_activation_function  is
	Port(
		neuron_output: in signed;
		activation_result
	);
end step_activation_function
